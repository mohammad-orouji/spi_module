library ieee;
use ieee.std_logic_1164.all;

entity top_tb is
end;

architecture testbench of top_tb is
       
signal enable_tb        : std_logic; 
signal reset_tb         : std_logic; 
signal clk_tb           : std_logic;
signal start_send_tb    : std_logic;
signal ERROR_TOP_tb     : std_logic_vector(3 downto 0);

constant T_10      : time    := 10    ns;

begin

    ins_0 : entity work.top
        port map(
            RESET_TOP       => reset_tb,
            CLK_TOP         => clk_tb,
            ENABLE_TOP      => enable_tb,
            START_SEN_TOP   => start_send_tb,
            ERROR_TOP       => ERROR_TOP_tb
        );

    process
    begin
        clk_tb  <= '0' ;
        wait for T_10/2;
        clk_tb  <= '1' ;
        wait for T_10/2;
    end process;

    reset_tb        <= '1'  , '0' after (T_10)/2, '1' after 20 us, '0' after 30 us ;
    enable_tb       <= '0'  , '1' after 50 ns;
    start_send_tb   <= '1' after 20 ns, '0' after 50 us;

end architecture testbench;